// 三速以太网MAC复位模块

module tri_mode_ethernet_mac_reset (


);

//------------------------------------
//             Local Signal
//------------------------------------


//------------------------------------
//             User Logic
//------------------------------------


//------------------------------------
//             Output Port
//------------------------------------



//------------------------------------
//             Instance
//------------------------------------


  endmodule