// PWM 参数配置模块, 解析参数并分发至相应通道
//   word 0: bit[ 7: 0] 通道索引
//           bit[31: 8] 保留
//   word 1: bit[31: 0] PWM输出频率, 单位Hz
//   word 2: bit[ 6: 0] PWM输出占空比, 0-100%
//           bit[31: 7] 保留
//   word 3: 保留
//   word 4: bit[ 0: 0] PWM输出使能
//           bit[31: 1] 保留

module pwm_config #(
  parameter   ID_PWM_PARAM = 0, // PWM参数帧ID
  parameter   CLK_FREQ = 100000000 // 模块时钟频率, Unit: Hz
)(
  // 模块时钟及复位
  input         clk,
  input         rst,
  // 用户UDP数据接收接口
  input  [31:0] rx_axis_udp_tdata,
  input         rx_axis_udp_tvalid,
  input         rx_axis_udp_tlast,
  input  [7:0]  rx_axis_udp_tuser, // 帧类型
  //输出参数
  output        pwm_config_vld, // 参数配置使能
  output [7:0]  pwm_config_channel, // 通道索引
  output        pwm_en, // PWM输出使能
  output [27:0] pwm_period, // 单周期计数时间
  output [27:0] pwm_hlevel // 高电平持续计数时间
);

//------------------------------------
//             Local Signal
//------------------------------------
  reg  [31:0]  rx_axis_udp_tdata_d1 = 0; // 打拍, 减小扇出
  reg          rx_axis_udp_tvalid_d1 = 0;
  reg          rx_axis_udp_tlast_d1 = 0;
  reg  [7:0]   word_cnt = 0; // word计数器
  reg          pwm_param_en = 0; // PWM参数帧使能
  reg  [27:0]  pwm_frequency = 0; // PWM输出频率
  reg  [6:0]   pwm_duty = 0; // PWM输出占空比
  reg          cal_period_en = 0; // 计算单周期计数时间使能
  reg          cal_period_en_d1 = 0; // 计算单周期计数时间使能
// 输出寄存器
  reg          pwm_config_vld_ff = 0; // 参数配置使能
  reg  [7:0]   pwm_config_channel_ff = 0; // 通道索引
  reg          pwm_en_ff = 0; // PWM输出使能
  reg  [27:0]  pwm_period_ff = 0; // 单周期计数时间
  reg  [27:0]  pwm_hlevel_ff = 0; // 高电平持续计数时间
//------------------------------------
//             User Logic
//------------------------------------
// 打拍, 减小扇出
  always @ (posedge clk) rx_axis_udp_tdata_d1 <= rx_axis_udp_tdata;
  always @ (posedge clk) rx_axis_udp_tvalid_d1 <= rx_axis_udp_tvalid;
  always @ (posedge clk) rx_axis_udp_tlast_d1 <= rx_axis_udp_tlast;

// 接收word计数器
  always @ (posedge clk)
    if (rst)
      word_cnt <= 0;
    else if (rx_axis_udp_tvalid_d1 && rx_axis_udp_tlast_d1)
      word_cnt <= 0;
    else if (rx_axis_udp_tvalid_d1)
      word_cnt <= word_cnt + 1; 
// 帧识别
  always @(posedge clk or posedge rst)
    if (rst)
      pwm_param_en <= 1'b0;
    else if (rx_axis_udp_tuser == ID_PWM_PARAM[7:0])
      pwm_param_en <= 1'b1;
    else
      pwm_param_en <= 1'b0;
// 参数解析
  // 通道索引
    always @ (posedge clk) if (pwm_param_en && (word_cnt == 0) && rx_axis_udp_tvalid_d1) pwm_config_channel_ff <= rx_axis_udp_tdata_d1[7:0];
  // PWM输出频率
    always @ (posedge clk) if (pwm_param_en && (word_cnt == 1) && rx_axis_udp_tvalid_d1) pwm_frequency <= rx_axis_udp_tdata_d1[27:0];
  // PWM输出占空比
    always @ (posedge clk) if (pwm_param_en && (word_cnt == 2) && rx_axis_udp_tvalid_d1) pwm_duty <= rx_axis_udp_tdata_d1[6:0];
  // PWM输出使能
    always @ (posedge clk) if (pwm_param_en && (word_cnt == 4) && rx_axis_udp_tvalid_d1) pwm_en_ff <= rx_axis_udp_tdata_d1[0];
// 计算单周期计数时间
  always @ (posedge clk)
    if (pwm_param_en && rx_axis_udp_tvalid_d1 && rx_axis_udp_tlast_d1)
      cal_period_en <= 1'b1;
    else if (m_axis_dout_tvalid)
      cal_period_en <= 1'b0;
  always @ (posedge clk) cal_period_en_d1 <= cal_period_en;

  always @ (posedge clk)
    if ((!cal_period_en_d1) && cal_period_en)
      begin
        s_axis_divisor_tvalid <= 1'b1;
        s_axis_divisor_tdata  <= {4'b0,pwm_frequency};
        s_axis_dividend_tvalid <= 1'b1;
        s_axis_dividend_tdata <= (CLK_FREQ[31:0] + {5'b0,pwm_frequency[27:1]}); // 四舍五入
      end
    else if (m_axis_dout_tvalid && cal_period_en)
      begin
        s_axis_divisor_tvalid <= 1'b1;
        s_axis_divisor_tdata  <= {4'b0,pwm_frequency};
        s_axis_dividend_tvalid <= 1'b1;
        s_axis_dividend_tdata <= ({5'b0,pwm_mul_p} + {6'b0,pwm_mul_p[26:1]}); // 四舍五入
      end
    else
      begin
        s_axis_divisor_tvalid <= 1'b0;
        s_axis_divisor_tdata  <= 32'b0;
        s_axis_dividend_tvalid <= 1'b0;
        s_axis_dividend_tdata <= 32'b0;
      end
  assign pwm_mul_a = pwm_duty;

//------------------------------------
//             Output Port
//------------------------------------
  assign pwm_config_vld     = pwm_config_vld;
  assign pwm_config_channel = pwm_config_channel;
  assign pwm_en             = pwm_en;
  assign pwm_period         = pwm_period;
  assign pwm_hlevel         = pwm_hlevel;

//------------------------------------
//             Instance
//------------------------------------
reg          s_axis_divisor_tvalid = 0;
reg  [31:0]  s_axis_divisor_tdata = 0;
reg          s_axis_dividend_tvalid = 0;
reg  [31:0]  s_axis_dividend_tdata = 0;
wire         m_axis_dout_tvalid;
wire [63:0]  m_axis_dout_tdata;
wire [6:0]   pwm_mul_a = 0;
wire [26:0]  pwm_mul_p = 0;
// Xilinx Divider Generate IP
  // Radix2, Unsigned 28bits / Unsigned 28bits, Remainder, Latency = 30 clocks
  div_gen_u28_u28 pwm_div(
    .aclk,
    // 除数
    .s_axis_divisor_tvalid,
    .s_axis_divisor_tdata,
    // 被除数
    .s_axis_dividend_tvalid,
    .s_axis_dividend_tdata,
    // 商+余数
    .m_axis_dout_tvalid,
    .m_axis_dout_tdata
  )
// Xilinx Multiplier IP
  mult_gen_x1000000 pwm_mul(
    .CLK(clk),
    .A  (pwm_mul_a),
    .P  (pwm_mul_p)
  )
  endmodule