// 三速以太网MAC复位模块

module pwm_ctrl (


);

//------------------------------------
//             Local Signal
//------------------------------------


//------------------------------------
//             User Logic
//------------------------------------


//------------------------------------
//             Output Port
//------------------------------------



//------------------------------------
//             Instance
//------------------------------------


  endmodule